`timescale 1ns/1ps

// TOP MODULE
module uart_top
#(
parameter clk_freq = 1000000,
parameter baud_rate = 9600
)
(
  input clk,rst, 
  input rx,
  input [7:0] dintx,
  input newd,
  output tx, 
  output [7:0] doutrx,
  output donetx,
  output donerx
    );
    
uarttx 
#(clk_freq, baud_rate) 
utx   
(clk, rst, newd, dintx, tx, donetx);   
 
uartrx 
#(clk_freq, baud_rate)
rtx
(clk, rst, rx, donerx, doutrx);    
    
endmodule
 

// TRANSMITTER MODULE
module uarttx
#(
    parameter clk_freq = 1000000 ,
    parameter baud_rate = 9600
)
(
    input clk, rst,
    input newd,
    input [7:0] tx_data,
    output reg tx,
    output reg donetx
);

localparam clkcount = clk_freq/baud_rate;
integer count=0;
integer counts=0;
reg uclk=0;

enum bit[1:0] {idle=2'b00, start=2'b01, transfer=2'b10, done=2'b11} state;

// UART clock generation
always @(posedge clk) begin
    if(count<clkcount/2) count<=count+1;
    else begin
        count=0;
        uclk<=~uclk;
    end
end

reg [7:0] din;

always @(posedge uclk) begin
    if(rst) state<=idle;
    else begin
        case (state)
        idle: begin
            counts<=0;
            tx<=1'b1;
            donetx<=1'b0;
            if(newd) begin
                state<=transfer;
                din<=tx_data;
                tx<=1'b0;
            end
            else state<=idle;
        end

        transfer: begin
            if(counts<=7) begin
                counts<=counts+1;
                tx<=din[counts];
                state<=transfer;
            end
            else begin
                counts<=0;
                tx<=1'b1;
                state<=idle;
                donetx<=1'b1;
            end
        end

        default: state<=idle;
        endcase
    end
end
endmodule

////////////////////

// RECIEVER MODULE
module uartrx
#(
    parameter clk_freq = 1000000 ,
    parameter baud_rate = 9600
)
(
    input clk, rst,
    input rx,
    output reg done,
    output reg [7:0] rxdata,
);

localparam clkcount = clk_freq/baud_rate;
integer count=0;
integer counts=0;
reg uclk=0;

enum bit[1:0] {idle=2'b00, start=2'b01} state;

// UART clock generation
always @(posedge clk) begin
    if(count<clkcount/2) count<=count+1;
    else begin
        count=0;
        uclk<=~uclk;
    end
end

always @(posedge uclk) begin
    if(rst)begin
        rxdata<=8'h00;
        counts<=0;
        done<=1'b0;
    end
    else begin
        case (state)
        idle: begin
            counts<=0;
            rxdata<=8'h00;
            done<=1'b0;
            if(rx==1'b0) begin
                state<=start;
            end
            else state<=idle;
        end

        start: begin
            if(counts<=7) begin
                counts<=counts+1;
                rxdata<={rx,rxdata[7:1]};
            end
            else begin
                counts<=0;
                done<=1'b1;
                state<=idle;
            end
        end

        default: state<=idle;
        endcase
    end
end
endmodule

///////////////////////////////////////////////////////////////////
 
interface uart_if;
  logic clk;
  logic uclktx;
  logic uclkrx;
  logic rst;
  logic rx;
  logic [7:0] dintx;
  logic newd;
  logic tx;
  logic [7:0] doutrx;
  logic donetx;
  logic donerx;
  
endinterface